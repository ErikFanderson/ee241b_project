VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_SPACING STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 4000 ;
END UNITS
MANUFACTURINGGRID 0.00025 ;

MACRO nem_sw
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN nem_sw 0 0 ;
  SIZE 0.096 BY 0.075 ;
  SYMMETRY X Y R90 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.038 0.057 0.056 0.075 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.038 0 0.056 0.018 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.078 0 0.096 0.018 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 0 0.018 0.018 ;
      LAYER M3 ;
        RECT 0 0 0.018 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.018 0.018 ;
      LAYER M1 ;
        RECT 0 0 0.018 0.018 ;
      LAYER V1 ;
        RECT 0 0 0.018 0.018 ;
      LAYER V2 ;
        RECT 0 0 0.018 0.018 ;
      LAYER V3 ;
        RECT 0 0 0.018 0.018 ;
    END
  END B
  OBS
    LAYER LIG SPACING 0.02 ;
      RECT 0 0 0.096 0.075 ;
    LAYER M1 SPACING 0.018 ;
      RECT 0 0.05 0.096 0.075 ;
      RECT 0.05 0 0.096 0.075 ;
    LAYER M2 SPACING 0.018 ;
      RECT 0 0.05 0.096 0.075 ;
      RECT 0.05 0 0.096 0.075 ;
    LAYER M3 ;
      RECT 0.078 0 0.096 0.075 ;
    LAYER M3 SPACING 0.018 ;
      RECT 0 0.05 0.096 0.075 ;
      RECT 0.05 0 0.096 0.075 ;
    LAYER M4 SPACING 0.018 ;
      RECT 0 0.05 0.096 0.075 ;
      RECT 0.05 0 0.096 0.075 ;
    LAYER M5 SPACING 0.018 ;
      RECT 0 0.05 0.096 0.075 ;
      RECT 0.05 0 0.096 0.075 ;
  END
END nem_sw

END LIBRARY
