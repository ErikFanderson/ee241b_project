//nems_sw.v
//DEPRECATED: REPLACED BY LEF

module nem_sw (
    inout wire [0:0] D,
    inout wire [0:0] S,
    input wire [0:0] G,
    input wire [0:0] B
    );

//define w/ lef


endmodule
