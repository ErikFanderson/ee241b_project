global vdd vss

.SUBCKT nem_sw D G S B 
r0 D net6 200 
r1 net6 S 200
c0 net6 vss 1e-13
.ENDS
