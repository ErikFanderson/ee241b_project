* SPICE NETLIST
***************************************

.SUBCKT nem_sw
** N=9 EP=0 IP=0 FDC=0
.ENDS
***************************************
