global vdd vss

.SUBCKT nem_sw D G S B 
r0 D net6 1e3
r1 net6 S 1e3
c0 net6 vss 1e-12
.ENDS
