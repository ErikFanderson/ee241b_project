.SUBCKT nems_relay drain gate source vss vdd
r0 drain net6 1e3
r1 net6 source 1e3
c0 net6 vss 1e-12
.ENDS
