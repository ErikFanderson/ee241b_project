VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_SPACING STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 4000 ;
END UNITS
MANUFACTURINGGRID 0.00025 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER well
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END well

LAYER Gate
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.02 ;
  AREA 0.06 ;
  SPACING 0.034 ;
  DIAGSPACING 0.19 ;
  PROPERTY LEF58_TYPE "TYPE POLYROUTING ;" ;
END Gate

LAYER Active
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
END Active

LAYER LISD
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE MEOL ;" ;
END LISD

LAYER LIG
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE MEOL ;" ;
END LIG

LAYER V0
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
END V0

LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 0.036 ;
  WIDTH 0.018 ;
  OFFSET 0.018 0.018 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0 0.018 ;
  MINIMUMCUT 1 WIDTH 0.01775 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMABOVE ;
  DIAGPITCH 0.051 0.051 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
END M1

LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.036 0.036 ;
  WIDTH 0.018 ;
  OFFSET 0.018 0.018 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0 0.018 ;
  MINIMUMCUT 1 WIDTH 0.01775 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMABOVE ;
  DIAGPITCH 0.051 0.051 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
END M2

LAYER V1
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
END V1

LAYER V2
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 0.036 ;
  WIDTH 0.018 ;
  OFFSET 0.018 0.018 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0 0.18 ;
  MINIMUMCUT 1 WIDTH 0.01775 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.01775 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMABOVE ;
  DIAGPITCH 0.051 0.051 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
END M3

LAYER V3
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.048 0.048 ;
  WIDTH 0.024 ;
  OFFSET 0.024 0.024 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0 0.024 ;
  MINIMUMCUT 1 WIDTH 0.01775 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.02375 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMABOVE ;
  DIAGPITCH 0.068 0.068 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
END M4

LAYER V4
  TYPE CUT ;
  SPACING 0.034 ;
  WIDTH 0.024 ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.048 0.048 ;
  WIDTH 0.024 ;
  OFFSET 0.024 0.024 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0 0.024 ;
  MINIMUMCUT 1 WIDTH 0.02375 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.02375 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMABOVE ;
  DIAGPITCH 0.068 0.068 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
END M5

LAYER V5
  TYPE CUT ;
  SPACING 0.034 ;
  WIDTH 0.024 ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.064 0.064 ;
  WIDTH 0.032 ;
  OFFSET 0.032 0.032 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0 0.032 ;
  MINIMUMCUT 1 WIDTH 0.02375 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.03175 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMABOVE ;
  DIAGPITCH 0.068 0.068 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
END M6

LAYER V6
  TYPE CUT ;
  SPACING 0.046 ;
  WIDTH 0.032 ;
END V6

LAYER M7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.064 0.064 ;
  WIDTH 0.032 ;
  OFFSET 0.032 0.032 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0 0.032 ;
  MINIMUMCUT 1 WIDTH 0.03175 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.12975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.13975 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.42475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1.14475 WITHIN 0.295 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.03175 WITHIN 1.705 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.35975 WITHIN 1.705 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.80475 WITHIN 1.705 FROMABOVE ;
  DIAGPITCH 0.068 0.068 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
END M7

LAYER V7
  TYPE CUT ;
  SPACING 0.046 ;
  WIDTH 0.032 ;
END V7

LAYER M8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 0.08 ;
  WIDTH 0.04 ;
  OFFSET 0.04 0.04 ;
  AREA 7.52 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.39975 1.19975 1.79975 
    WIDTH 0 0.04 0.04 0.04 0.04 
    WIDTH 0.05975 0.04 0.06 0.04 0.04 
    WIDTH 0.07975 0.04 0.04 0.08 0.04 
    WIDTH 0.11975 0.04 0.04 0.04 0.12 
    WIDTH 0.49975 0.04 0.04 0.04 0.5 
    WIDTH 0.99975 0.04 0.04 0.04 1 ;
  MINIMUMCUT 1 WIDTH 0.03175 WITHIN 1.705 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.35975 WITHIN 1.705 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.80475 WITHIN 1.705 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.03975 WITHIN 1.705 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.35975 WITHIN 1.705 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.80475 WITHIN 1.705 FROMABOVE ;
  MAXWIDTH 2 ;
  MINSTEP 0.04 STEP ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 20 20 ;
  DENSITYCHECKSTEP 10 ;
END M8

LAYER V8
  TYPE CUT ;
  SPACING 0.057 ;
  WIDTH 0.04 ;
END V8

LAYER SDT
  TYPE CUT ;
END SDT

LAYER M9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.08 0.08 ;
  WIDTH 0.04 ;
  OFFSET 0.04 0.04 ;
  AREA 7.52 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.39975 1.19975 1.79975 
    WIDTH 0 0.04 0.04 0.04 0.04 
    WIDTH 0.05975 0.04 0.06 0.04 0.04 
    WIDTH 0.07975 0.04 0.04 0.08 0.04 
    WIDTH 0.11975 0.04 0.04 0.04 0.12 
    WIDTH 0.49975 0.04 0.04 0.04 0.5 
    WIDTH 0.99975 0.04 0.04 0.04 1 ;
  MINIMUMCUT 1 WIDTH 0.03975 WITHIN 1.705 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0.35975 WITHIN 1.705 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.80475 WITHIN 1.705 FROMABOVE ;
  MAXWIDTH 2 ;
  MINSTEP 0.04 STEP ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 80 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M9

LAYER V9
  TYPE CUT ;
  SPACING 0.057 ;
  WIDTH 0.04 ;
END V9

LAYER Pad
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 0.08 ;
  WIDTH 0.04 ;
  OFFSET 0.04 0.04 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 11.99975 
    WIDTH 0 2 2 
    WIDTH 11.99975 2 3 ;
  MINIMUMCUT 1 WIDTH 0.03975 WITHIN 1.705 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.35975 WITHIN 1.705 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.80475 WITHIN 1.705 FROMBELOW ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 80 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END Pad

VIARULE Pad_M9 GENERATE DEFAULT
  LAYER M9 ;
    ENCLOSURE 0 0.011 ;
  LAYER Pad ;
    ENCLOSURE 0.011 0 ;
  LAYER V9 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.078 BY 0.078 ;
END Pad_M9

VIARULE M9_M8 GENERATE DEFAULT
  LAYER M8 ;
    ENCLOSURE 0.02 0 ;
  LAYER M9 ;
    ENCLOSURE 0 0.02 ;
  LAYER V8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
    SPACING 0.097 BY 0.097 ;
END M9_M8

VIARULE M8_M7 GENERATE DEFAULT
  LAYER M7 ;
    ENCLOSURE 0 0.011 ;
  LAYER M8 ;
    ENCLOSURE 0.011 0 ;
  LAYER V7 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.078 BY 0.078 ;
END M8_M7

VIARULE M7_M6 GENERATE DEFAULT
  LAYER M6 ;
    ENCLOSURE 0.011 0 ;
  LAYER M7 ;
    ENCLOSURE 0 0.011 ;
  LAYER V6 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.078 BY 0.078 ;
END M7_M6

VIARULE M6_M5 GENERATE DEFAULT
  LAYER M5 ;
    ENCLOSURE 0 0.011 ;
  LAYER M6 ;
    ENCLOSURE 0.011 0 ;
  LAYER V5 ;
    RECT -0.012 -0.012 0.012 0.012 ;
    SPACING 0.058 BY 0.058 ;
END M6_M5

VIARULE M5_M4 GENERATE DEFAULT
  LAYER M4 ;
    ENCLOSURE 0.011 0 ;
  LAYER M5 ;
    ENCLOSURE 0 0.011 ;
  LAYER V4 ;
    RECT -0.012 -0.012 0.012 0.012 ;
    SPACING 0.058 BY 0.058 ;
END M5_M4

VIARULE M4_M3 GENERATE DEFAULT
  LAYER M3 ;
    ENCLOSURE 0 0.005 ;
  LAYER M4 ;
    ENCLOSURE 0.011 0 ;
  LAYER V3 ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.036 BY 0.036 ;
END M4_M3

VIARULE M3_M2 GENERATE DEFAULT
  LAYER M2 ;
    ENCLOSURE 0.005 0 ;
  LAYER M3 ;
    ENCLOSURE 0 0.005 ;
  LAYER V2 ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.036 BY 0.036 ;
END M3_M2

VIARULE M2_M1 GENERATE DEFAULT
  LAYER M1 ;
    ENCLOSURE 0 0.005 ;
  LAYER M2 ;
    ENCLOSURE 0.005 0 ;
  LAYER V1 ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.036 BY 0.036 ;
END M2_M1

SITE coreSite
  CLASS CORE ;
  SYMMETRY X R90 ;
  SIZE 0.054 BY 0.27 ;
END coreSite

MACRO nem_sw
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN nem_sw 0 0 ;
  SIZE 0.096 BY 0.075 ;
  SYMMETRY X Y R90 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.038 0.057 0.056 0.075 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.038 0 0.056 0.018 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.078 0 0.096 0.018 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0 0 0.018 0.018 ;
      LAYER M3 ;
        RECT 0 0 0.018 0.018 ;
      LAYER M2 ;
        RECT 0 0 0.018 0.018 ;
      LAYER M1 ;
        RECT 0 0 0.018 0.018 ;
      LAYER V1 ;
        RECT 0 0 0.018 0.018 ;
      LAYER V2 ;
        RECT 0 0 0.018 0.018 ;
      LAYER V3 ;
        RECT 0 0 0.018 0.018 ;
    END
  END B
  OBS
    LAYER LIG SPACING 0.02 ;
      RECT 0 0 0.096 0.075 ;
    LAYER M1 SPACING 0.018 ;
      RECT 0 0.05 0.096 0.075 ;
      RECT 0.05 0 0.096 0.075 ;
    LAYER M2 SPACING 0.018 ;
      RECT 0 0.05 0.096 0.075 ;
      RECT 0.05 0 0.096 0.075 ;
    LAYER M3 ;
      RECT 0.078 0 0.096 0.075 ;
    LAYER M3 SPACING 0.018 ;
      RECT 0 0.05 0.096 0.075 ;
      RECT 0.05 0 0.096 0.075 ;
  END
END nem_sw

END LIBRARY
